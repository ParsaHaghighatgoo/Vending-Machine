`timescale 1ns / 1ps

module supportphase(
    );

initial begin
str1="you can send ur opinin to us or what u want with send an email to example@gmail.com";
$display("str1 = %s",str1);

endmodule
